version https://git-lfs.github.com/spec/v1
oid sha256:26cde97e3259e22b7ca0a6624c92eaf8f099efa216d7dd7dc6a7989514c6520f
size 5111
