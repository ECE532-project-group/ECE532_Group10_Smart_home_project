version https://git-lfs.github.com/spec/v1
oid sha256:12b7684e02c6562f74b31154ec84852285b308922035f6444889d5ec3bf5e2ae
size 11689
