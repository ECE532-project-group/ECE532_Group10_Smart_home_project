version https://git-lfs.github.com/spec/v1
oid sha256:e6b8c5983dad9142df834f806db9294551218b2cc92964be906c6f3a2e2003b1
size 5567
