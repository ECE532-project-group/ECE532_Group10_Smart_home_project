version https://git-lfs.github.com/spec/v1
oid sha256:4c16c11ab37300180f7dbe41da75f41627cbebd1110aa694962f6fa1f6ce67ca
size 5827
