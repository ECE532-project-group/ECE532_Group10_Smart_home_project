version https://git-lfs.github.com/spec/v1
oid sha256:729d371150b3a69fe183fb5fd50121a4129a6377b930708917a93ef20cf8a217
size 4872
